`define L2_ASSOCIATIVITY 2
`define L2_SETS 8
`define L2_W_INDEX $clog2(`L2_SETS)

`define D_ASSOCIATIVITY 4
`define D_SETS 8
`define D_W_INDEX $clog2(`D_SETS)

`define I_ASSOCIATIVITY 4
`define I_SETS 8
`define I_W_INDEX $clog2(`I_SETS)